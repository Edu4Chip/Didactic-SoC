`INCREMENT_CYCLE_COUNT(clk_i)
