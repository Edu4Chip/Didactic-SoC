`INCREMENT_CYCLE_COUNT(clk_in)
`include "verification/verilator/src/generated/hdl/ms/Student_SS_3_0.sv"
