`INCREMENT_CYCLE_COUNT(clk)
`include "verification/verilator/src/generated/hdl/ms/Student_SS_2_0.sv"
