//-----------------------------------------------------------------------------
// File          : SS_Ctrl_reg_array.v
// Creation date : 23.02.2024
// Creation time : 12:38:00
// Description   :
// Created by    :
// Tool : Kactus2 3.13.1 64-bit
// Plugin : Verilog generator 2.4
// This file was generated based on IP-XACT component tuni.fi:ip:SS_Ctrl_reg_array:1.0
// whose XML file is C:/Users/kayra/Documents/repos/tau-ipxact/ipxact/tuni.fi/ip/SS_Ctrl_reg_array/1.0/SS_Ctrl_reg_array.1.0.xml
//-----------------------------------------------------------------------------
/*
  Contributors:
    * Matti Käyrä (matti.kayra@tuni.fi)
  Description:
    * Interface generated by kactus2, then manually continued and edited
    * This initial created manually.
    * same functionality can be later created by TAU Kamel tool automatically from IPXACT
*/


module SS_Ctrl_reg_array #(
    parameter IOCELL_CFG_W     = 5,
    parameter IOCELL_COUNT     = 28, // update/propagate this value to match cell numbers
    parameter AW = 32,
    parameter DW = 32,
    parameter SS_CTRL_W = 31, // configurable up to 31 bits
    parameter NUM_SS = 4
) (

    // Interface: Clock
    input  logic clk,

    // Interface: Reset
    input  logic reset_n,

    // Interface: icn_ss_ctrl
    output logic [SS_CTRL_W-1:0] ss_ctrl_icn,

    // Interface: io_cfg
    output logic [(IOCELL_CFG_W*IOCELL_COUNT)-1:0] cell_cfg,

    // Interface: mem_reg_if
    input  logic [AW-1:0]   addr_i,
    input  logic [DW/8-1:0] be_i,
    input  logic            req_i,
    input  logic [DW-1:0]   wdata_i,
    input  logic            we_i,
    input  logic            rready_i,
    output logic [DW-1:0]   rdata_o,
    output logic            rvalid_o,
    output logic            rvalidpar_o,
    output logic            gnt_o,
    output logic            gntpar_o,

    // Interface: rst_icn
    output logic reset_icn,

    // Interface: rst_ss_0
    output logic [NUM_SS-1:0] reset_ss,

    // Interface: ss_ctrl_0
    output logic                 irq_en_0,
    output logic [SS_CTRL_W-1:0] ss_ctrl_0,

    // Interface: ss_ctrl_1
    output logic                 irq_en_1,
    output logic [SS_CTRL_W-1:0] ss_ctrl_1,

    // Interface: ss_ctrl_2
    output logic                 irq_en_2,
    output logic [SS_CTRL_W-1:0] ss_ctrl_2,

    // Interface: ss_ctrl_3
    output logic                 irq_en_3,
    output logic [SS_CTRL_W-1:0] ss_ctrl_3,

    // Interface: ss_ctrl_4
    output logic                 irq_en_4,
    output logic [SS_CTRL_W-1:0] ss_ctrl_4,

    // Interface: pmod_ctrl
    output logic [7:0] pmod_sel,

    // Interface: fetch_en
    output logic [3:0] fetch_en
);


  logic [31:0] fetch_en_reg;
  logic [31:0] ss_rst_reg;
  logic [31:0] icn_ctrl_reg;
  logic [31:0] ss_0_ctrl_reg;
  logic [31:0] ss_1_ctrl_reg;
  logic [31:0] ss_2_ctrl_reg;
  logic [31:0] ss_3_ctrl_reg;
  logic [31:0] ss_4_ctrl_reg;
  logic [31:0] ss_ctrl_reserved_1_reg;
  logic [31:0] pmod_sel_reg;
  // gpio layout: uart/spi/gpio
  logic [IOCELL_COUNT-1:0][31:0] io_cell_cfg_reg;

  logic [31:0] boot_reg_0;
  logic [31:0] boot_reg_1;
  logic [31:0] return_reg_0;
  logic [31:0] return_reg_1;

  logic rvalid_reg;
  logic gnt_reg;
  logic [DW-1:0] rdata_out_reg;

    // FFs for write or read/write registers
    always_ff @( posedge clk or negedge reset_n )
    begin : control_register_ff
    if (~reset_n) begin
        fetch_en_reg <= 'h5;
        ss_rst_reg <= 'h0;
        icn_ctrl_reg <= 'h0;
        ss_0_ctrl_reg <= 'h0;
        ss_1_ctrl_reg <= 'h0;
        ss_2_ctrl_reg <= 'h0;
        ss_3_ctrl_reg <= 'h0;
        ss_4_ctrl_reg <= 'h0;
        ss_ctrl_reserved_1_reg <= 'h0;
        pmod_sel_reg <= 'h4;
        for(int i=0; i < IOCELL_COUNT; i++) begin
          io_cell_cfg_reg[i] <= 'h0;
        end
        boot_reg_0 <= 'h6f;
        boot_reg_1 <= 'h6f;
        return_reg_0 <= 'h6f;
        return_reg_1 <= 'h6f;

        rvalid_reg <= 1'b0;
        gnt_reg <= 1'b1;
        rdata_out_reg <= 'h0;
        
    end
    else begin

      // req - gnt handshake
      if(req_i & gnt_reg) begin
        gnt_reg <= 1'b0;
      end

      if (we_i & req_i & ~rvalid_reg) begin

        // io cell cfg
        for(int i=0; i < IOCELL_COUNT; i++) begin
          if ( addr_i == 'h28+i*4) begin // check 28 - 88
            io_cell_cfg_reg[i] <= wdata_i;
          end
        end

        case (addr_i[16:0])
          'h0:  fetch_en_reg <= wdata_i;
          'h4:  ss_rst_reg   <= wdata_i;

          'h8:  icn_ctrl_reg           <= wdata_i;
          'hC:  ss_0_ctrl_reg          <= wdata_i;
          'h10: ss_1_ctrl_reg          <= wdata_i;
          'h14: ss_2_ctrl_reg          <= wdata_i;
          'h18: ss_3_ctrl_reg          <= wdata_i;
          'h1C: ss_4_ctrl_reg          <= wdata_i;

          'h20: ss_ctrl_reserved_1_reg <= wdata_i;

          'h24: pmod_sel_reg <= wdata_i;

          //unrolled io cells conf would be here

          'h100: boot_reg_0   <= wdata_i;
          'h104: boot_reg_1   <= wdata_i;
          'h180: return_reg_0 <= wdata_i;
          'h184: return_reg_1 <= wdata_i;
        endcase

        rvalid_reg <= 1'b1;
      end
      else if(~we_i & req_i & ~rvalid_reg) begin 

        for(int i=0; i < IOCELL_COUNT; i++) begin
          if ( addr_i == 'h28+i*4) begin // check 28 - 88
              rdata_out_reg <= io_cell_cfg_reg[i];
          end
        end

        // io cell cfg
        case(addr_i[16:0])

          'h0:  rdata_out_reg <= fetch_en_reg;
          'h4:  rdata_out_reg <= ss_rst_reg;

          'h8:  rdata_out_reg <= icn_ctrl_reg;
          'hC:  rdata_out_reg <= ss_0_ctrl_reg;
          'h10: rdata_out_reg <= ss_1_ctrl_reg;
          'h14: rdata_out_reg <= ss_2_ctrl_reg;
          'h18: rdata_out_reg <= ss_3_ctrl_reg;
          'h1C: rdata_out_reg <= ss_4_ctrl_reg;

          'h20: rdata_out_reg <= ss_ctrl_reserved_1_reg;

          'h24: rdata_out_reg <= pmod_sel_reg;

          //unrolled io cells conf would be here

          'h100: rdata_out_reg <= boot_reg_0;
          'h104: rdata_out_reg <= boot_reg_1;
          'h180: rdata_out_reg <= return_reg_0;
          'h184: rdata_out_reg <= return_reg_1;
 
        endcase
        rvalid_reg <= 1'b1;
      end
      else if(~rready_i & ~gnt_reg) begin
        rvalid_reg <= 1'b1;
      end
      else begin
        gnt_reg    <= 1'b1;
        rvalid_reg <= 1'b0;
      end
    end
  end // control_register_ff

  always_comb // 
  begin : comb_logic
    
    rvalid_o    = rvalid_reg;
    rvalidpar_o = ~rvalid_reg;
    gnt_o       = gnt_reg;
    gntpar_o    = ~gnt_reg;
    rdata_o     = rdata_out_reg;

    for(int i=0; i < IOCELL_COUNT; i++) begin
      cell_cfg[i*IOCELL_CFG_W +:IOCELL_CFG_W] = io_cell_cfg_reg[i];
    end

end // comb_logic

// assign ins - potential status regs that can be read

// assign outs

assign reset_icn  = ss_rst_reg[0];
assign reset_ss = ss_rst_reg[NUM_SS:1];

assign irq_en_0    = ss_0_ctrl_reg[31];
assign ss_ctrl_0   = ss_0_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_1    = ss_1_ctrl_reg[31];
assign ss_ctrl_1   = ss_1_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_2    = ss_2_ctrl_reg[31] ;
assign ss_ctrl_2   = ss_2_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_3    = ss_3_ctrl_reg[31];
assign ss_ctrl_3   = ss_3_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_4    = ss_4_ctrl_reg[31];
assign ss_ctrl_4   = ss_4_ctrl_reg[SS_CTRL_W-1:0];
assign ss_ctrl_icn = icn_ctrl_reg[SS_CTRL_W-1:0];

assign pmod_sel = pmod_sel_reg;

assign fetch_en = fetch_en_reg[3:0];

// this functionality can be recreated by kamel framework once memory design is finalized.
// ipxact register map needs to be synced to this rtl first
endmodule
