`INCREMENT_CYCLE_COUNT(clk)
`include "verification/verilator/src/generated/hdl/ms/SysCtrl_peripherals_0.sv"
