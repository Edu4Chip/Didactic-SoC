`INCREMENT_CYCLE_COUNT(clk_i)
`include "verification/verilator/src/generated/hdl/ms/jtag_dbg_wrapper.sv"
