`include "verification/verilator/src/common.v"
`INCREMENT_CYCLE_COUNT(clk_i)
