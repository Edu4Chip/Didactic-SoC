`INCREMENT_CYCLE_COUNT(clk)
`include "verification/verilator/src/generated/hdl/ms/AX4LITE_APB_converter_wrapper.sv"
