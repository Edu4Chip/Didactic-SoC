`INCREMENT_CYCLE_COUNT(clock)
