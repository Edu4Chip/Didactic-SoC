`INCREMENT_CYCLE_COUNT(clk)
