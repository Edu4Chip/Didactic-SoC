`INCREMENT_CYCLE_COUNT(clock)
`include "verification/verilator/src/generated/hdl/ms/SysCtrl_SS_wrapper_0.sv"
