module VipDidactic #()();
endmodule : VipDidactic
