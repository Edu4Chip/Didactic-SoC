`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/Student_SS_1_0.sv"
