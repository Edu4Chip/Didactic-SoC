`INCREMENT_CYCLE_COUNT(clk_i)
`include "verification/verilator/src/generated/hdl/ms/mem_axi_bridge.sv"
