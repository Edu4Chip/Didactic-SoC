`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/student_ss_1.sv"
