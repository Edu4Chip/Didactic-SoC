//-----------------------------------------------------------------------------
// File          : ICN_SS.v
// Creation date : 19.02.2024
// Creation time : 15:01:06
// Description   : 
// Created by    : 
// Tool : Kactus2 3.13.1 64-bit
// Plugin : Verilog generator 2.4
// This file was generated based on IP-XACT component tuni.fi:interconnect:ICN_SS:1.0
// whose XML file is C:/Users/kayra/Documents/repos/tau-ipxact/ipxact/tuni.fi/interconnect/ICN_SS/1.0/ICN_SS.1.0.xml
//-----------------------------------------------------------------------------
/*
  Contributors:
    * Matti Käyrä (matti.kayra@tuni.fi)
  Description:
    * example "interconnect"
    * interface generated by kactus2
*/
module ICN_SS #(
    parameter                              APB_AW           = 32,
    parameter                              APB_DW           = 32,
    parameter                              APB_TARGETS      = 4,
    parameter                              AXI_AW           = 32,
    parameter                              AXI_DW           = 32,
    parameter                              AXI_IDW          = 10,
    parameter                              AXI_USERW        = 1
) (
    // Interface: AXI
    input                [AXI_AW-1:0]   AR_ADDR,
    input                [1:0]          AR_BURST,
    input                [3:0]          AR_CACHE,
    input                [AXI_IDW-1:0]  AR_ID,
    input                [7:0]          AR_LEN,
    input                               AR_LOCK,
    input                [2:0]          AR_PROT,
    input                [3:0]          AR_QOS,
    input                [2:0]          AR_REGION,
    input                [2:0]          AR_SIZE,
    input                [AXI_USERW-1:0] AR_USER,
    input                               AR_VALID,
    input                [AXI_AW-1:0]   AW_ADDR,
    input                [5:0]          AW_ATOP,
    input                [1:0]          AW_BURST,
    input                [3:0]          AW_CACHE,
    input                [AXI_IDW-1:0]  AW_ID,
    input                [7:0]          AW_LEN,
    input                               AW_LOCK,
    input                [2:0]          AW_PROT,
    input                [3:0]          AW_QOS,
    input                [3:0]          AW_REGION,
    input                [2:0]          AW_SIZE,
    input                [AXI_USERW-1:0] AW_USER,
    input                               AW_VALID,
    input                               B_READY,
    input                               R_READY,
    input                [AXI_DW-1:0]   W_DATA,
    input                               W_LAST,
    input                [(AXI_DW/8)-1:0] W_STROBE,
    input                [AXI_USERW-1:0] W_USER,
    input                               W_VALID,
    output                              AR_READY,
    output                              AW_READY,
    output               [AXI_IDW-1:0]  B_ID,
    output               [1:0]          B_RESP,
    output               [AXI_USERW-1:0] B_USER,
    output                              B_VALID,
    output               [AXI_DW-1:0]   R_DATA,
    output               [AXI_IDW-1:0]  R_ID,
    output                              R_LAST,
    output               [1:0]          R_RESP,
    output               [AXI_USERW-1:0] R_USER,
    output                              R_VALID,
    output                              W_READY,

    // Interface: Clock
    input                               clk,

    // Interface: Reset
    input                               reset_int,

    // Interface: SS_Ctrl
    input                [7:0]          ss_ctrl_icn,

    // There ports are contained in many interfaces
    input                [(APB_DW*APB_TARGETS)-1:0] PRDATA,
    input                [APB_TARGETS-1:0] PREADY,
    input                [APB_TARGETS-1:0] PSLVERR,
    output               [APB_AW-1:0]   PADDR,
    output                              PENABLE,
    output               [APB_TARGETS-1:0] PSEL,
    output               [APB_DW-1:0]   PWDATA,
    output                              PWRITE
);

  // TODO: FIll parameters
  AXI_BUS #(
    .AXI_ADDR_WIDTH(), 
    .AXI_DATA_WIDTH(), 
    .AXI_ID_WIDTH(), 
    .AXI_USER_WIDTH()
  ) axi4bus ();

  AXI_LITE #(
   .AXI_ADDR_WIDTH(),
   .AXI_DATA_WIDTH()
  ) axi4lite_bus ();

  axi_to_axi_lite_intf #(

  )
  i_axi_to_axi_lite(
    .clk_i(clk),
    .rst_ni(reset_int),
    .testmode_i(1'b0),
    .slv(axi4bus),
    .mst(axi4lite_bus)
  );

  // TODO: Assign axi to interface
  assign axi4bus.ar_addr = AR_ADDR;





  //  APB addr decoding
  localparam APB_TARGETS=4;
  localparam NoAddrRules =4;
  localparam ADDR_BASE=32'h1300_0000
  localparam APB_SIZE='h1000;

  typedef axi_pkg::xbar_rule_32_t rule_t;

  rule_t [NoAddrRules-1:0] AddrMapAPB;
  // TODO: finalize Address table based on APB Subsystems
  assign AddrMapAPB = '{
                         '{idx: 32'd3, start_addr: ADDR_BASE+APB_SIZE*3, end_addr: ADDR_BASE+APB_SIZE*4-1},
                         '{idx: 32'd2, start_addr: ADDR_BASE+APB_SIZE*2, end_addr: ADDR_BASE+APB_SIZE*3-1},
                         '{idx: 32'd1, start_addr: ADDR_BASE+APB_SIZE*1, end_addr: ADDR_BASE+APB_SIZE*2-1},
                         '{idx: 32'd0, start_addr: ADDR_BASE+APB_SIZE*0, end_addr: ADDR_BASE+APB_SIZE*1-1}
                         };

  // TODO: fill parameters
  axi_lite_to_apb_intf #(
    .NoApbSlaves(),
    .NoRules(),
    .AddrWidth(),
    .DataWidth(),
    .rule_t(rule_t)
    )
  i_axi_lite_to_apb_intf(
    .clk_i(clk),
    .rst_ni(reset_int),

    .slv(axi4lite_bus),

    .paddr_o(PADDR),
    .pprot_o(),
    .pselx_o(PSEL),
    .penable_o(PENABLE),
    .pwrite_o(PWRITE),
    .pwdata_o(PWDATA),
    .pstrb_o(),
    .pready_i(PREADY),
    .prdata_i(PRDATA),
    .pslverr_i(PSLVERR),

    .addr_map_i(AddrMapAPB)
  );


endmodule
