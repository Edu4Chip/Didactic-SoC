`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/SS_Ctrl_reg_array.sv"
