//-----------------------------------------------------------------------------
// File          : io_cell_frame_ss_1.v
// Creation date : 15.02.2024
// Creation time : 15:30:39
// Description   : 
// Created by    : 
// Tool : Kactus2 3.13.1 64-bit
// Plugin : Verilog generator 2.4
// This file was generated based on IP-XACT component tuni.fi:subsystem.io:io_cell_frame_ss_1:1.0
// whose XML file is C:/Users/kayra/Documents/repos/tau-ipxact/tuni.fi/subsystem.io/io_cell_frame_ss_1/1.0/io_cell_frame_ss_1.1.0.xml
//-----------------------------------------------------------------------------

module io_cell_frame_ss_1(
    // Interface: GPIO_external
    inout                [1:0]          gpio,

    // Interface: GPIO_internal
    input                [1:0]          gpio_oe,
    input                [1:0]          gpo_in,
    output               [1:0]          gpi_out,

    // These ports are not in any interface
    input                [4:0]          io_cell_cfg
);

// WARNING: EVERYTHING ON AND ABOVE THIS LINE MAY BE OVERWRITTEN BY KACTUS2!!!
endmodule
