`include "verification/verilator/src/generated/hdl/ms/pmod_mux.sv"
