`INCREMENT_CYCLE_COUNT(clk)
`include "verification/verilator/src/generated/hdl/ms/Student_SS_0_0.sv"
