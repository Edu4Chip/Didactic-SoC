`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/AX4LITE_APB_converter_wrapper.sv"
