`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/SysCtrl_xbar.sv"
