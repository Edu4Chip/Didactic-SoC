`INCREMENT_CYCLE_COUNT(clk)
`include "verification/verilator/src/generated/hdl/ms/ICN_SS.sv"
