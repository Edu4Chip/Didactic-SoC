`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/jtag_dbg_wrapper.sv"
