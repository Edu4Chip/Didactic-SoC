`INCREMENT_CYCLE_COUNT(clk_internal)
`include "verification/verilator/src/generated/hdl/ms/SysCtrl_SS_0.sv"
