`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/ibex_axi_bridge.sv"
