//-----------------------------------------------------------------------------
// File          : SS_Ctrl_reg_array.v
// Creation date : 23.02.2024
// Creation time : 12:38:00
// Description   :
// Created by    :
// Tool : Kactus2 3.13.1 64-bit
// Plugin : Verilog generator 2.4
// This file was generated based on IP-XACT component tuni.fi:ip:SS_Ctrl_reg_array:1.0
// whose XML file is C:/Users/kayra/Documents/repos/tau-ipxact/ipxact/tuni.fi/ip/SS_Ctrl_reg_array/1.0/SS_Ctrl_reg_array.1.0.xml
//-----------------------------------------------------------------------------
/*
  Contributors:
    * Matti Käyrä (matti.kayra@tuni.fi)
  Description:
    * Interface generated by kactus2, then manually continued and edited
    * This initial created manually.
    * same functionality can be later created by TAU Kamel tool automatically from IPXACT
*/


module SS_Ctrl_reg_array #(
    parameter IOCELL_CFG_W     = 5,
    parameter IOCELL_COUNT     = 28, // update/propagate this value to match cell numbers
    parameter AW = 32,
    parameter DW = 32,
    parameter SS_CTRL_W = 31 // configurable up to 31 bits
) (

    // Interface: Clock
    input  logic clk,

    // Interface: Reset
    input  logic reset,

    // Interface: icn_ss_ctrl
    output logic [SS_CTRL_W-1:0]          ss_ctrl_icn,

    // Interface: io_cfg
    output logic [(IOCELL_CFG_W*IOCELL_COUNT)-1:0] cell_cfg,

    // Interface: mem_reg_if
    input  logic [AW-1:0]   addr_in,
    input  logic [DW/8-1:0] be_in,
    input  logic            req_in,
    input  logic [DW-1:0]   wdata_in,
    input  logic            we_in,
    output logic [DW-1:0]   rdata_out,

    // Interface: rst_icn
    output logic reset_icn,

    // Interface: rst_ss_0
    output logic reset_ss_0,

    // Interface: rst_ss_1
    output logic reset_ss_1,

    // Interface: rst_ss_2
    output logic reset_ss_2,

    // Interface: rst_ss_3
    output logic reset_ss_3,

    // Interface: ss_ctrl_0
    output logic                 irq_en_0,
    output logic [SS_CTRL_W-1:0] ss_ctrl_0,

    // Interface: ss_ctrl_1
    output logic                 irq_en_1,
    output logic [SS_CTRL_W-1:0] ss_ctrl_1,

    // Interface: ss_ctrl_2
    output logic                 irq_en_2,
    output logic [SS_CTRL_W-1:0] ss_ctrl_2,

    // Interface: ss_ctrl_3
    output logic                 irq_en_3,
    output logic [SS_CTRL_W-1:0] ss_ctrl_3,

    // Interface: pmod_ctrl
    output logic [7:0] pmod_sel,

    // Interface: fetch_en
    output logic [4:0] fetch_en
);


  logic [31:0] fetch_en_reg;
  logic [31:0] ss_rst_reg;
  logic [31:0] icn_ctrl_reg;
  logic [31:0] ss_0_ctrl_reg;
  logic [31:0] ss_1_ctrl_reg;
  logic [31:0] ss_2_ctrl_reg;
  logic [31:0] ss_3_ctrl_reg;
  logic [31:0] ss_ctrl_reserved_0_reg;
  logic [31:0] ss_ctrl_reserved_1_reg;
  logic [31:0] pmod_sel_reg;
  logic [IOCELL_COUNT-1:0][31:0] io_cell_cfg_reg;

  logic [31:0] boot_reg_0;
  logic [31:0] boot_reg_1;
  logic [31:0] return_reg_0;
  logic [31:0] return_reg_1;

    // FFs for write or read/write registers
    always_ff @( posedge clk or negedge reset )
    begin : control_register_ff
    if (~reset) begin
        fetch_en_reg <= 'h5;
        ss_rst_reg <= 'h0;
        icn_ctrl_reg <= 'h0;
        ss_0_ctrl_reg <= 'h0;
        ss_1_ctrl_reg <= 'h0;
        ss_2_ctrl_reg <= 'h0;
        ss_3_ctrl_reg <= 'h0;
        ss_ctrl_reserved_0_reg <= 'h0;
        ss_ctrl_reserved_1_reg <= 'h0;
        pmod_sel_reg <= 'h4;
        for(int i=0; i < IOCELL_COUNT; i++) begin
          io_cell_cfg_reg[i] <= 'h0;
        end
        boot_reg_0 <= 'h6f;
        boot_reg_1 <= 'h6f;
        return_reg_0 <= 'h6f;
        return_reg_1 <= 'h6f;
    end
    else begin

     if (we_in) begin
        case (addr_in[16:0])
        'h0:  fetch_en_reg       <= wdata_in;
        'h4:  ss_rst_reg         <= wdata_in;

        'h8:  icn_ctrl_reg       <= wdata_in;
        'hC:  ss_0_ctrl_reg      <= wdata_in;
        'h10: ss_1_ctrl_reg      <= wdata_in;
        'h14: ss_2_ctrl_reg      <= wdata_in;
        'h18: ss_3_ctrl_reg      <= wdata_in;

        'h1C: ss_ctrl_reserved_0_reg <= wdata_in;
        'h20: ss_ctrl_reserved_1_reg <= wdata_in;

        'h24: pmod_sel_reg        <= wdata_in;

        'h28: io_cell_cfg_reg[0]  <= wdata_in;
        'h2C: io_cell_cfg_reg[1]  <= wdata_in;
        'h30: io_cell_cfg_reg[2]  <= wdata_in;
        'h34: io_cell_cfg_reg[3]  <= wdata_in;

        'h38: io_cell_cfg_reg[4]  <= wdata_in;
        'h3C: io_cell_cfg_reg[5]  <= wdata_in;
        'h40: io_cell_cfg_reg[6]  <= wdata_in;
        'h44: io_cell_cfg_reg[7]  <= wdata_in;

        'h48: io_cell_cfg_reg[8]  <= wdata_in;
        'h4C: io_cell_cfg_reg[9]  <= wdata_in;
        'h50: io_cell_cfg_reg[10] <= wdata_in;
        'h54: io_cell_cfg_reg[11] <= wdata_in;
        'h58: io_cell_cfg_reg[12] <= wdata_in;
        'h5C: io_cell_cfg_reg[13] <= wdata_in;
        'h60: io_cell_cfg_reg[14] <= wdata_in;

        'h64: io_cell_cfg_reg[15] <= wdata_in;
        'h68: io_cell_cfg_reg[16] <= wdata_in;

        //'h6C: io_cell_cfg_reg[17] <= wdata_in;
        //'h70: io_cell_cfg_reg[18] <= wdata_in;

        'h100: boot_reg_0 <= wdata_in;
        'h104: boot_reg_1 <= wdata_in;
        'h180: return_reg_0 <= wdata_in;
        'h184: return_reg_1 <= wdata_in;

        endcase
     end
    end
    end // control_register_ff

    always_comb // read process
    begin : read_logic
      rdata_out = 'h0;
      case(addr_in[16:0])

        'h0:  rdata_out = fetch_en_reg;
        'h4:  rdata_out = ss_rst_reg;

        'h8:  rdata_out = icn_ctrl_reg;
        'hC:  rdata_out = ss_0_ctrl_reg;
        'h10: rdata_out = ss_1_ctrl_reg;
        'h14: rdata_out = ss_2_ctrl_reg;
        'h18: rdata_out = ss_3_ctrl_reg;

        'h1C: rdata_out = ss_ctrl_reserved_0_reg;
        'h20: rdata_out = ss_ctrl_reserved_1_reg;

        'h24: rdata_out = pmod_sel_reg;
        // gpio 0
        'h28: rdata_out = io_cell_cfg_reg[0];
        'h2C: rdata_out = io_cell_cfg_reg[1];
        'h30: rdata_out = io_cell_cfg_reg[2];
        'h34: rdata_out = io_cell_cfg_reg[3];
        // gpio 1
        'h38: rdata_out = io_cell_cfg_reg[4];
        'h3C: rdata_out = io_cell_cfg_reg[5];
        'h40: rdata_out = io_cell_cfg_reg[6];
        'h44: rdata_out = io_cell_cfg_reg[7];
        // spi
        'h48: rdata_out = io_cell_cfg_reg[8];
        'h4C: rdata_out = io_cell_cfg_reg[9];
        'h50: rdata_out = io_cell_cfg_reg[10];
        'h54: rdata_out = io_cell_cfg_reg[11];
        'h58: rdata_out = io_cell_cfg_reg[12];
        'h5C: rdata_out = io_cell_cfg_reg[13];
        'h60: rdata_out = io_cell_cfg_reg[14];
        // uart
        'h64: rdata_out = io_cell_cfg_reg[15];
        'h68: rdata_out = io_cell_cfg_reg[16];
        // reserves
        //'h6C: rdata_out = io_cell_cfg_reg[17];
        //'h70: rdata_out = io_cell_cfg_reg[18];

        'h100: rdata_out = boot_reg_0;
        'h104: rdata_out = boot_reg_1;
        'h180: rdata_out = return_reg_0;
        'h184: rdata_out = return_reg_1;

    endcase

    for(int i=0; i < IOCELL_COUNT; i++) begin
      cell_cfg[i*IOCELL_CFG_W +:IOCELL_CFG_W] = io_cell_cfg_reg[i];
    end
end // read_logic

// assign ins


// assign outs

assign reset_icn  = ss_rst_reg[0];
assign reset_ss_0 = ss_rst_reg[1];
assign reset_ss_1 = ss_rst_reg[2];
assign reset_ss_2 = ss_rst_reg[3];
assign reset_ss_3 = ss_rst_reg[4];

assign irq_en_0    = ss_0_ctrl_reg[31];
assign ss_ctrl_0   = ss_0_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_1    = ss_1_ctrl_reg[31];
assign ss_ctrl_1   = ss_1_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_2    = ss_2_ctrl_reg[31] ;
assign ss_ctrl_2   = ss_2_ctrl_reg[SS_CTRL_W-1:0];
assign irq_en_3    = ss_3_ctrl_reg[31];
assign ss_ctrl_3   = ss_3_ctrl_reg[SS_CTRL_W-1:0];
assign ss_ctrl_icn = icn_ctrl_reg[SS_CTRL_W-1:0];

assign pmod_sel = pmod_sel_reg;

assign fetch_en = fetch_en_reg[4:0];

// this functionality can be recreated by kamel framework once memory design is finalized.
// ipxact register map needs to be synced to this rtl first
endmodule
