`include "verification/verilator/src/common.v"
