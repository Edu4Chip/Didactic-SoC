`INCREMENT_CYCLE_COUNT(clk_in)
