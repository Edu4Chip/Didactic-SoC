`include "verification/verilator/src/hdl/common.v"
`include "verification/verilator/src/generated/hdl/nms/Student_area_0.sv"
