//-----------------------------------------------------------------------------
// File          : jtag_dbg_wrapper.v
// Creation date : 16.02.2024
// Creation time : 12:34:42
// Description   : 
// Created by    : 
// Tool : Kactus2 3.13.1 64-bit
// Plugin : Verilog generator 2.4
// Interface was originally generated based on IP-XACT component tuni.fi:ip:jtag_dbg_wrapper:1.0
//-----------------------------------------------------------------------------
/*
  Contributors:
    * Antti Nurmi    (antti.nurmi@tuni.fi)
    * Tom Szymkowiak (thomas.szymkowiak@tuni.fi)
    * Matti Käyrä    (matti.kayra@tuni.fi)
  Description:
    * debug module intergration wrapper
    * interface generated by kactus2
    * original module implementation by AN and TZS
    * tweaks for importing to kactus2 by MK
*/

module jtag_dbg_wrapper #(
    parameter                              AXI_AW           = 32,
    parameter                              AXI_DW           = 32,
    parameter                              DM_BASE_ADDRESS  = 'h1000,
    parameter                              DM_ID_VALUE  =  32'hf007ba11
  )(
    // Interface: AXI4LITE_I
    input  logic                  init_ar_ready,
    input  logic                  init_aw_ready,
    input  logic [1:0]            init_b_resp,
    input  logic                  init_b_valid,
    input  logic [AXI_DW-1:0]     init_r_data,
    input  logic [1:0]            init_r_resp,
    input  logic                  init_r_valid,
    input  logic                  init_w_ready,
    output logic [AXI_AW-1:0]     init_ar_addr,
    output logic                  init_ar_valid,
    output logic [3:0]            init_ar_prot,
    output logic [AXI_AW-1:0]     init_aw_addr,
    output logic                  init_aw_valid,
    output logic [3:0]            init_aw_prot,
    output logic                  init_b_ready,
    output logic                  init_r_ready,
    output logic [AXI_DW-1:0]     init_w_data,
    output logic [(AXI_DW/8)-1:0] init_w_strb,
    output logic                  init_w_valid,

    // Interface: AXI4LITE_T
    input  logic [AXI_AW-1:0]     target_ar_addr,
    input  logic                  target_ar_valid,
    input  logic [AXI_AW-1:0]     target_aw_addr,
    input  logic                  target_aw_valid,
    input  logic                  target_b_ready,
    input  logic                  target_r_ready,
    input  logic [AXI_DW-1:0]     target_w_data,
    input  logic [(AXI_DW/8)-1:0] target_w_strb,
    input  logic                  target_w_valid,
    output logic                  target_ar_ready,
    output logic                  target_aw_ready,
    output logic [1:0]            target_b_resp,
    output logic                  target_b_valid,
    output logic [AXI_DW-1:0]     target_r_data,
    output logic [1:0]            target_r_resp,
    output logic                  target_r_valid,
    output logic                  target_w_ready,

    // Interface: Clock
    input  logic                  clk_i,

    // Interface: Debug
    output logic                  debug_req_irq_o,

    // Interface: JTAG
    input  logic                  jtag_tck_i,
    input  logic                  jtag_td_i,
    input  logic                  jtag_tms_i,
    input  logic                  jtag_trst_ni,
    output logic                  jtag_td_o,

    // Interface: Reset
    input  logic                  rstn_i,

    // Interface: core_reset
    output logic                  core_reset,

    // These ports are not in any interface
    output logic                  ndmreset_o
  );

/****** LOCAL VARIABLES AND CONSTANTS *****************************************/

localparam int unsigned NrHarts       =  1;
localparam int unsigned DBG_BUS_WIDTH = 32;

// static debug hartinfo
localparam dm::hartinfo_t DebugHartInfo = '{
  zero1:                 '0,
  nscratch:               2, // Debug module needs at least two scratch regs
  zero0:                 '0,
  dataaccess:          1'b1, // data registers are memory mapped in the debugger
  datasize:   dm::DataCount,
  dataaddr:   dm::DataAddr
};

// JTAG TAP <-> DMI signals
dm::dmi_req_t                 dmi_req_s;
dm::dmi_resp_t                dmi_resp_s;
logic                         dmi_req_valid_s;
logic                         dmi_req_ready_s;
logic                         dmi_resp_valid_s;
logic                         dmi_resp_ready_s;
// dbg_s 
logic                         dbg_s_req_s;
logic                         dbg_s_we_s;
logic [DBG_BUS_WIDTH-1:0]     dbg_s_addr_s;
logic [DBG_BUS_WIDTH-1:0]     dbg_s_wdata_s;
logic [(DBG_BUS_WIDTH/8)-1:0] dbg_s_be_s;
logic [DBG_BUS_WIDTH-1:0]     dbg_s_rdata_s;
// dbg_m
logic                         dbg_m_req_s;
logic [DBG_BUS_WIDTH-1:0]     dbg_m_add_s;
logic                         dbg_m_we_s;
logic [DBG_BUS_WIDTH-1:0]     dbg_m_wdata_s;
logic [DBG_BUS_WIDTH/8-1:0]   dbg_m_be_s;
logic                         dbg_m_gnt_s;
logic                         dbg_m_valid_s;
logic [DBG_BUS_WIDTH-1:0]     dbg_m_rdata_s;

/****** COMPONENT + INTERFACE INSTANTIATIONS **********************************/

  ibex_axi_bridge #(
    .AXI_AW ( AXI_AW ),
    .AXI_DW ( AXI_DW ),
    .IBEX_AW( DBG_BUS_WIDTH  ),
    .IBEX_DW( DBG_BUS_WIDTH  )
  ) i_debug2axi_lite_bridge (
    .clk_i      ( clk_i                   ),
    .rst_ni     ( rstn_i                  ),
    .req_i      ( dbg_m_req_s             ),
    .gnt_o      ( dbg_m_gnt_s             ),
    .rvalid_o   ( dbg_m_valid_s           ),
    .we_i       ( dbg_m_we_s              ),
    .be_i       ( dbg_m_be_s              ),
    .addr_i     ( dbg_m_add_s             ),
    .wdata_i    ( dbg_m_wdata_s           ),
    .rdata_o    ( dbg_m_rdata_s           ),
    .err_o      ( /* NC */                ),
    .aw_addr_o  ( init_aw_addr  ),
    .aw_valid_o ( init_aw_valid ),
    .aw_ready_i ( init_aw_ready ),
    .w_data_o   ( init_w_data   ),
    .w_strb_o   ( init_w_strb   ),
    .w_valid_o  ( init_w_valid  ),
    .w_ready_i  ( init_w_ready  ),
    .b_resp_i   ( init_b_resp   ),
    .b_valid_i  ( init_b_valid  ),
    .b_ready_o  ( init_b_ready  ),
    .ar_addr_o  ( init_ar_addr  ),
    .ar_valid_o ( init_ar_valid ),
    .ar_ready_i ( init_ar_ready ),
    .r_data_i   ( init_r_data   ),
    .r_resp_i   ( init_r_resp   ),
    .r_valid_i  ( init_r_valid  ),
    .r_ready_o  ( init_r_ready  )
  );

  assign init_aw_prot = '0;
  assign init_ar_prot = '0;

  mem_axi_bridge #(
    .MEM_AW    ( DBG_BUS_WIDTH ),
    .MEM_DW    ( DBG_BUS_WIDTH ),
    .AXI_AW    ( AXI_AW        ),
    .AXI_DW    ( AXI_DW        ),
    .ADDR_MASK ( 'h0           )
  ) i_axi_lite2debug_bridge (
    .clk_i      ( clk_i             ),
    .rst_ni     ( rstn_i            ),
    .req_o      ( dbg_s_req_s       ),
    .we_o       ( dbg_s_we_s        ),
    .addr_o     ( dbg_s_addr_s      ),
    .wdata_o    ( dbg_s_wdata_s     ),
    .be_o       ( dbg_s_be_s        ),
    .rdata_i    ( dbg_s_rdata_s     ),
    .aw_addr_i  ( target_aw_addr    ),
    .aw_valid_i ( target_aw_valid   ),
    .aw_ready_o ( target_aw_ready   ),
    .w_data_i   ( target_w_data     ),
    .w_strb_i   ( target_w_strb     ),
    .w_valid_i  ( target_w_valid    ),
    .w_ready_o  ( target_w_ready    ),
    .b_resp_o   ( target_b_resp     ),
    .b_valid_o  ( target_b_valid    ),
    .b_ready_i  ( target_b_ready    ),
    .ar_addr_i  ( target_ar_addr    ),
    .ar_valid_i ( target_ar_valid   ),
    .ar_ready_o ( target_ar_ready   ),
    .r_data_o   ( target_r_data     ),
    .r_resp_o   ( target_r_resp     ),
    .r_valid_o  ( target_r_valid    ),
    .r_ready_i  ( target_r_ready    )
  );


  dmi_jtag #(
    .IdcodeValue (DM_ID_VALUE)
  ) i_dmi_jtag (
    .clk_i                ( clk_i            ),
    .rst_ni               ( rstn_i           ),
    .testmode_i           ( '0               ),
    .dmi_rst_no           ( /*nc*/           ),
    .dmi_req_valid_o      ( dmi_req_valid_s  ),
    .dmi_req_ready_i      ( dmi_req_ready_s  ),
    .dmi_req_o            ( dmi_req_s        ),
    .dmi_resp_valid_i     ( dmi_resp_valid_s ),
    .dmi_resp_ready_o     ( dmi_resp_ready_s ),
    .dmi_resp_i           ( dmi_resp_s       ),
    .tck_i                ( jtag_tck_i       ),
    .tms_i                ( jtag_tms_i       ),
    .trst_ni              ( jtag_trst_ni     ),
    .td_i                 ( jtag_td_i        ),
    .td_o                 ( jtag_td_o        ),
    .tdo_oe_o             ( /*nc*/           )
  );

  dm_top #(
    .NrHarts         ( NrHarts         ),  
    .BusWidth        ( DBG_BUS_WIDTH   ),   
    .DmBaseAddress   ( DM_BASE_ADDRESS ), // TBD     
    .SelectableHarts ( {NrHarts{1'b1}} ),          
    .ReadByteEnable  ( 1               ) // toggle new behavior to drive master_be_o during a read    
  ) i_dm_top (
    .clk_i                ( clk_i               ),
    .rst_ni               ( rstn_i              ),
    .testmode_i           ( '0                  ),
    .ndmreset_o           ( ndmreset_o          ),
    .ndmreset_ack_i       ( '0                  ),//new feature of dm_top
    .dmactive_o           ( /*nc*/              ),
    .debug_req_o          ( debug_req_irq_o     ),
    .unavailable_i        ( '0                  ),
    .hartinfo_i           ( DebugHartInfo       ),
    .slave_req_i          ( dbg_s_req_s         ),
    .slave_we_i           ( dbg_s_we_s          ),
    .slave_addr_i         ( dbg_s_addr_s        ),
    .slave_be_i           ( dbg_s_be_s          ),
    .slave_wdata_i        ( dbg_s_wdata_s       ),
    .slave_rdata_o        ( dbg_s_rdata_s       ),
    .master_req_o         ( dbg_m_req_s         ),
    .master_add_o         ( dbg_m_add_s         ),
    .master_we_o          ( dbg_m_we_s          ),
    .master_wdata_o       ( dbg_m_wdata_s       ),
    .master_be_o          ( dbg_m_be_s          ),
    .master_gnt_i         ( dbg_m_gnt_s         ),
    .master_r_valid_i     ( dbg_m_valid_s       ),
    .master_r_rdata_i     ( dbg_m_rdata_s       ),
    .master_r_other_err_i ( '0                  ),
    .master_r_err_i       ( '0                  ),
    .dmi_rst_ni           ( rstn_i              ),
    .dmi_req_valid_i      ( dmi_req_valid_s     ),
    .dmi_req_ready_o      ( dmi_req_ready_s     ),
    .dmi_req_i            ( dmi_req_s           ),
    .dmi_resp_valid_o     ( dmi_resp_valid_s    ),
    .dmi_resp_ready_i     ( dmi_resp_ready_s    ),
    .dmi_resp_o           ( dmi_resp_s          )
  );

  // ibex core reset control with debug module
  assign core_reset = rstn_i & ~(ndmreset_o);

endmodule
